module color_control(hcounter, vcounter, mouse_x, mouse_y, map, val_red, val_green, val_blue);

input [9:0] hcounter, vcounter, mouse_x, mouse_y;
input [5:0] map [99:0];
output reg [3:0] val_red, val_green, val_blue;

reg [63:0] block_empty [47:0];
reg [63:0] block_bomb [47:0];
reg [63:0] block_1 [47:0];
reg [63:0] block_2 [47:0];
reg [63:0] block_3 [47:0];
reg [63:0] block_4 [47:0];

reg [1:0] color;    // 0: white, 1: black, 2: grey;
wire [3:0] row_coor, col_coor;
wire i_val, j_val;

assign col_coor = (hcounter - 144) / 64;
assign row_coor = (vcounter - 35) / 48;
assign j_val = (hcounter - 144) % 64;
assign i_val = (vcounter - 35) % 48;

initial begin
    block_empty = '{
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111
    };
    block_bomb = '{
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000011111100000000000000000000001111,
        64'b1111000000000000000000000000001111111111000000000110000000001111,
        64'b1111000000000000000000000000011110001111100000001110000000001111,
        64'b1111000000000000000000000000111100000011110000001110000000001111,
        64'b1111000000000000000000000000111000000001111000011100000000001111,
        64'b1111000000000000000000000001111000000000111111111000000000001111,
        64'b1111000000000000000000000111111110000000001111110000000000001111,
        64'b1111000000000000000000111111111111110000000000000000000000001111,
        64'b1111000000000000000001111100000011111000000000000000000000001111,
        64'b1111000000000000000011100000000000011100000000000000000000001111,
        64'b1111000000000000000111000000000000001110000000000000000000001111,
        64'b1111000000000000001110000000000000000111000000000000000000001111,
        64'b1111000000000000011100000000000000000011100000000000000000001111,
        64'b1111000000000000111000000000000000000001110000000000000000001111,
        64'b1111000000000000110000000000000000000000110000000000000000001111,
        64'b1111000000000000110000000000000000000000110000000000000000001111,
        64'b1111000000000001110000000000000000000000111000000000000000001111,
        64'b1111000000000001100000000000000000000000011000000000000000001111,
        64'b1111000000000001100000000000000000000000011000000000000000001111,
        64'b1111000000000001100000000000000000000000011000000000000000001111,
        64'b1111000000000001100000000000000000000000011000000000000000001111,
        64'b1111000000000001100000000000000000000000011000000000000000001111,
        64'b1111000000000001100000000000000000000000011000000000000000001111,
        64'b1111000000000001110000000000000000000000111000000000000000001111,
        64'b1111000000000000110000000000000000000000110000000000000000001111,
        64'b1111000000000000110000000000000000000000110000000000000000001111,
        64'b1111000000000000111000000000000000000001110000000000000000001111,
        64'b1111000000000000011100000000000000000011100000000000000000001111,
        64'b1111000000000000001110000000000000000111000000000000000000001111,
        64'b1111000000000000000111000000000000001110000000000000000000001111,
        64'b1111000000000000000011100000000000011100000000000000000000001111,
        64'b1111000000000000000001111100000011111000000000000000000000001111,
        64'b1111000000000000000000111111111111110000000000000000000000001111,
        64'b1111000000000000000000000111111110000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111
    };
    block_1 = '{
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111
    };
    block_2 = '{
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000000000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111
    };
    block_3 = '{
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000001111111111100000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111
    };
    block_4 = '{
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000111100000000000011110000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000011111111111100000000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000011110000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111000000000000000000000000000000000000000000000000000000001111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111,
        64'b1111111111111111111111111111111111111111111111111111111111111111
    };
end

always @(*) begin
    if(col_coor >= 10 || col_coor >= 10) begin
        color <= 2;
    end
    else begin
        case(map[row_coor * 10 + col_coor]) 
            6'b010001: color <= block_1[i][j];
            6'b010010: color <= block_2[i][j];
            6'b010011: color <= block_3[i][j];
            6'b010100: color <= block_4[i][j];
            6'b011000: color <= block_bomb[i][j];
            6'b110001: color <= block_empty[i][j];
            6'b110010: color <= block_empty[i][j];
            6'b110011: color <= block_empty[i][j];
            default: begin
                color = (0 <= i_val && i_val <= 3) || (44 <= i_val && i_val <= 47) || (0 <= j_val && j_val <= 3) || (60 <= j_val && j_val <= 63) ? 1 : 2;
            end
        endcase
    end
end

always @(*) begin
    case(color) 
        2'b00: begin
            val_red <= 4'b0000;
            val_green <= 4'b0000;
            val_blue <= 4'b0000;
        end
        2'b01: begin
            val_red <= 4'b1111;
            val_green <= 4'b1111;
            val_blue <= 4'b1111;
        end
        default: begin
            val_red <= 4'b0101;
            val_green <= 4'b0101;
            val_blue <= 4'b0101;
        end
    endcase
end

endmodule